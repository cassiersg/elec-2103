
module qsys1 (
	clk_clk,
	mtl_touch_ip_0_mtl_connection_i2cclock,
	mtl_touch_ip_0_mtl_connection_interruptic,
	mtl_touch_ip_0_mtl_connection_i2cdata,
	reset_reset_n);	

	input		clk_clk;
	output		mtl_touch_ip_0_mtl_connection_i2cclock;
	input		mtl_touch_ip_0_mtl_connection_interruptic;
	inout		mtl_touch_ip_0_mtl_connection_i2cdata;
	input		reset_reset_n;
endmodule
